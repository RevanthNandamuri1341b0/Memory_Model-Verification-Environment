/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 06 August 2021
*Time of update : 13:44
*Project name : MEMORY DUT VERIFICATION
*Domain : UVM
*Description : 
File Name : sequencer.sv
*File ID : 689645
*Modified by : #your name#
*/

typedef uvm_sequencer #(packet) sequencer;
