/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 04 October 2021
*Project name : Verification of Memory Model using RAL Verification
*Domain : UVM
*Description : 
*File Name : sequencer.sv
*File ID : 836883
*Modified by : #your name#
*/

typedef uvm_sequencer #(packet) sequencer;
