/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 05 October 2021
*Project name : Verification of Memory Model using RAL Verification with Backdoor access
*Domain : UVM
*Description : 
*File Name : sequencer.sv
*File ID : 336224
*Modified by : #your name#
*/

typedef uvm_sequencer #(packet) sequencer;